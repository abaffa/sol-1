library verilog;
use verilog.vl_types.all;
entity microcode_sequencer_sv_unit is
end microcode_sequencer_sv_unit;
