package pa_cpu;
  
  parameter PAGETABLE_RAM_SIZE = 2 ** 13;


endpackage
