library verilog;
use verilog.vl_types.all;
entity pa_microcode is
end pa_microcode;
