library verilog;
use verilog.vl_types.all;
entity pa_testbench is
end pa_testbench;
