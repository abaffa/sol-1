library verilog;
use verilog.vl_types.all;
entity pa_cpu is
end pa_cpu;
