library verilog;
use verilog.vl_types.all;
entity cpu_top_sv_unit is
end cpu_top_sv_unit;
