library verilog;
use verilog.vl_types.all;
entity microcode_sequencer is
    port(
        arst            : in     vl_logic;
        clk             : in     vl_logic;
        ir              : in     vl_logic_vector(7 downto 0);
        alu_flags       : in     vl_logic_vector(7 downto 0);
        cpu_status      : in     vl_logic_vector(7 downto 0);
        alu_out         : in     vl_logic_vector(7 downto 0);
        z_bus           : in     vl_logic_vector(7 downto 0);
        alu_of          : in     vl_logic;
        alu_final_cf    : in     vl_logic;
        dma_req         : in     vl_logic;
        \WAIT\          : in     vl_logic;
        int_pending     : in     vl_logic;
        ext_input       : in     vl_logic;
        u_flags         : out    vl_logic_vector(7 downto 0);
        ctrl_typ        : out    vl_logic_vector(1 downto 0);
        ctrl_offset     : out    vl_logic_vector(6 downto 0);
        ctrl_cond_invert: out    vl_logic;
        ctrl_cond_flag_src: out    vl_logic;
        ctrl_cond_sel   : out    vl_logic_vector(3 downto 0);
        ctrl_escape     : out    vl_logic;
        ctrl_u_zf_in_src: out    vl_logic_vector(1 downto 0);
        ctrl_u_cf_in_src: out    vl_logic_vector(1 downto 0);
        ctrl_u_sf_in_src: out    vl_logic;
        ctrl_u_of_in_src: out    vl_logic;
        ctrl_ir_wrt     : out    vl_logic;
        ctrl_status_flags_wrt: out    vl_logic;
        ctrl_shift_msb_src: out    vl_logic_vector(2 downto 0);
        ctrl_zbus_in_src_0: out    vl_logic_vector(1 downto 0);
        ctrl_alu_a_src  : out    vl_logic_vector(5 downto 0);
        ctrl_alu_op     : out    vl_logic_vector(3 downto 0);
        ctrl_alu_mode   : out    vl_logic;
        ctrl_alu_cf_in_src: out    vl_logic_vector(1 downto 0);
        ctrl_alu_cf_in_invert: out    vl_logic;
        ctrl_alu_cf_out_invert: out    vl_logic;
        ctrl_zf_in_src  : out    vl_logic_vector(1 downto 0);
        ctrl_cf_in_src  : out    vl_logic_vector(2 downto 0);
        ctrl_sf_in_src  : out    vl_logic_vector(1 downto 0);
        ctrl_of_in_src  : out    vl_logic_vector(2 downto 0);
        ctrl_rd         : out    vl_logic;
        ctrl_wr         : out    vl_logic;
        ctrl_alu_b_src  : out    vl_logic_vector(2 downto 0);
        ctrl_display_reg_load: out    vl_logic;
        ctrl_dl_wrt     : out    vl_logic;
        ctrl_dh_wrt     : out    vl_logic;
        ctrl_cl_wrt     : out    vl_logic;
        ctrl_ch_wrt     : out    vl_logic;
        ctrl_bl_wrt     : out    vl_logic;
        ctrl_bh_wrt     : out    vl_logic;
        ctrl_al_wrt     : out    vl_logic;
        ctrl_ah_wrt     : out    vl_logic;
        ctrl_mdr_in_src : out    vl_logic;
        ctrl_mdr_out_src: out    vl_logic;
        ctrl_mdr_out_en : out    vl_logic;
        ctrl_mdr_l_wrt  : out    vl_logic;
        ctrl_mdr_h_wrt  : out    vl_logic;
        ctrl_tdr_l_wrt  : out    vl_logic;
        ctrl_tdr_h_wrt  : out    vl_logic;
        ctrl_di_l_wrt   : out    vl_logic;
        ctrl_di_h_wrt   : out    vl_logic;
        ctrl_si_l_wrt   : out    vl_logic;
        ctrl_si_h_wrt   : out    vl_logic;
        ctrl_mar_l_wrt  : out    vl_logic;
        ctrl_mar_h_wrt  : out    vl_logic;
        ctrl_bp_l_wrt   : out    vl_logic;
        ctrl_bp_h_wrt   : out    vl_logic;
        ctrl_pc_l_wrt   : out    vl_logic;
        ctrl_pc_h_wrt   : out    vl_logic;
        ctrl_sp_l_wrt   : out    vl_logic;
        ctrl_sp_h_wrt   : out    vl_logic;
        ctrl_gl_wrt     : out    vl_logic;
        ctrl_gh_wrt     : out    vl_logic;
        ctrl_int_vector_wrt: out    vl_logic;
        ctrl_mask_flags_wrt: out    vl_logic;
        ctrl_mar_in_src : out    vl_logic;
        ctrl_int_ack    : out    vl_logic;
        ctrl_clear_all_ints: out    vl_logic;
        ctrl_ptb_wrt    : out    vl_logic;
        ctrl_page_table_we: out    vl_logic;
        ctrl_mdr_to_pagetable_data_buffer: out    vl_logic;
        ctrl_force_user_ptb: out    vl_logic;
        ctrl_immy       : out    vl_logic_vector(7 downto 0)
    );
end microcode_sequencer;
